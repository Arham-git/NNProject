module hello (
input a,
input b,
output c
);

c <= b + a;

endmodule